--
-- VHDL Entity ProjectWasmachine.test.arch_name
--
-- Created:
--          by - Perij.UNKNOWN (LAPTOP-Q0P13GKH)
--          at - 12:00:36 05/02/2025
--
-- using Mentor Graphics HDL Designer(TM) 2022.1 Built on 21 Jan 2022 at 13:00:30
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY test IS
END ENTITY test;

